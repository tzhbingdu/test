module test
(
input a,
output b
);

assign b=a;
assign c=a;

endmodule